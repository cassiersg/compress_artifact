`include "design.vh"
