module aes_round_umsk
(
    input [127:0] state,
    input [127:0] key,
    output 
);

endmodule
